module ysyx_22050243_ALUCTRL (
    input     
    input
    output reg [3:0] alu_ctrl
);