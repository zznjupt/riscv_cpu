module ysyx_22050243_id (
    input  wire             clk,
    input  wire             rst,
    input  wire [5:0]       stall,
    output wire             

);