module ysyx_22050243_REGSLICE # (
    parameter DATA_WIDTH = 1
) (
    input clk,
    input rst,
    
)